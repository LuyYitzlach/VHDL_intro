--this is the median sort shell
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.array_setup.all;


entity median_sort_VHDL is
generic (
	   numSize : integer := 33;
	   buffSize : integer := 6
		); --omit in tb
port 	(
		inBuff : in buffArray(numSize-1 downto 0)(buffSize-1 downto 0);
		clock  : in std_logic;
		outBuff : out buffArray(numSize-1 downto 0)(buffSize-1 downto 0);
		median : out std_logic_vector (numSize-1 downto 0)
		); --separate by ; but no ; on last item in () –omit in tb
end median_sort_VHDL;

architecture arch of median_sort_VHDL is
--declarations (type, signal, record, constants, components)
signal ii,jj,kk : integer;
--signal j : integer;
signal temp : std_logic_vector(numSize-1 downto 0);
signal temp_array : buffArray(numSize-1 downto 0)(buffSize-1 downto 0); 
constant half : integer := buffSize/2;

--procedures and functions
begin
process
begin 
-- procedure sorting (
		-- signal toSortArray : in buffArray(numSize-1 downto 0)(buffSize-1 downto 0);
		-- signal sortedArray : out buffArray(numSize-1 downto 0)(buffSize-1 downto 0)
		-- ) is
--signals for use within procedure

--begin
--put instructions for procedure here
 

	for k in 3 downto 1 loop --for k  in  half downto 1 loop
	kk <= k;
		for i  in 0 to 33 loop --for i  in 0 to buffSize loop
			ii <= i;
			jj <= ii+kk;
			if (jj < buffSize-1) then
				if (temp_array(ii) > temp_array(jj)) then
				temp <= temp_array(ii);
				wait for 10 ns; --add?
				temp_array(ii) <= temp_array(jj);
				temp_array(jj) <= temp; --how does this work if it's synchronous?
				--temp_array(i) <= temp_array(j);
				--temp_array(j) <= temp_array(i);
				end if;
			end if;
		ii <= ii+1;
		end loop;
	kk <= kk-1;
	exit when (kk = 0);
	end loop;
	
	
--sortedArray = temp_array;
--end sorting; --procedure ends
end process;

--processes, with their (local) variables
--instantiation/components (these could also be in declaration section)
--combinatorial expressions
temp_array <= inBuff;
--sorting(toSortArray => inBuff, sortedArray => outBuff);
median <= outBuff(2); --should really use division and flooring to find middle...
end arch;
